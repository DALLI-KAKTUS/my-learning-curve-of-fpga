`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    01:52:34 02/19/2023 
// Design Name: 
// Module Name:    inputs 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module inputs(
    input [3:0] switches_in,
	 output [3:0] switches_out
    );
	assign switches_in = switches_out;

endmodule
